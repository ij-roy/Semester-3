Hello IJ Roy