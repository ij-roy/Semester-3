Hello IJ